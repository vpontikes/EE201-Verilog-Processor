// Program memory implemented as combinational logic
// On the iCE40, this will be implemented in the logic fabric

// This is only used for the single-cycle machine; once we move to the
// multi-cycle design we will have a unified (and clocked) memory.

module progmem(input logic[31:0] addr,
               output logic[31:0] instr);

    // In the future, we will implement this by reading instructions stored in
    // an external file (which could be generated by an assembler), but for now
    // just hard-code the instructions here.
    // You can use Ripes to generate the bytes for the instructions you'd like
    // to run.

    // Code explanation:
    // 6 mod 4 (2) goes into x1, which is then subtracted from 10 (in x2), answ of 8 stored in x1

    always_comb
      case(addr)
        32'h0:  instr = 32'h00600093; // li x1, 6
        32'h4:  instr = 32'h00a00113; // li x2, 10
        32'h8:  instr = 32'h0030f093; // andi x1, x1, 0b11
        32'hc:  instr = 32'h401100b3; // sub x1, x2, x1
      default: instr = 0;
    endcase

endmodule

